
interface serializer_if;
    logic send_data_valid;
    logic [SEND_DATA_WIDTH-1:0] v_data_read;

endinterface
